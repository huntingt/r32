interface RVPair;
    logic ready;
    logic valid;


endinterface
